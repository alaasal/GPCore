package main;
    import uvm_package::*;
    `include "uvm_macros.svh"

    import pkg_memory::*;

    `include"core-component/c_core_agent_config.svh"
    `include"core-component/c_core_driver.svh"
    `include"core-component/c_core_request.svh"
    `include"core-component/c_core_monitor.svh"
    `include"core-component/c_core_agent.svh"
    `include"core-component/c_core_env.svh"
    `include"core-component/c_core_test.svh"
endpackage