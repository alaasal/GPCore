class memory_write_transaction extends memory_transaction;
   `uvm_object_utils(memory_write_transaction)

    t_write_op write_op;
    
endclass : memory_write_transaction
