package main;
    import uvm_package::*;
    `include "uvm_macros.svh"
    
endpackage