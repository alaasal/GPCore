class memory_read_transaction extends memory_transaction;
   `uvm_object_utils(memory_read_transaction)
;
    t_read_op read_op;
    
endclass : memory_read_transaction
