import pkg_memory::*;
import uvm_pkg::*;
`include"uvm_macros.svh"

module top ();
  
  initial begin
    run_test("memory_test");
  end
  
endmodule
