package main;
    import uvm_package::*;
    `include "uvm_macros.svh"

    import pkg_memory::*;

    `include"c_core_agent_config.svh"
    `include"c_core_driver.svh"
    `include"c_core_request.svh"
    `include"c_core_monitor.svh"
    `include"c_core_agent.svh"
endpackage